///////////////////////////////////////////////////////////////////////////////////
//																			     //
//  Copyright 2015-2016 by YanSolutions											 //
//                                                                               //
//  All rights reserved. The source code contained herein is publicly released   //
//  under the terms and conditions of the YanSolutions License. No part of       //
//  this source code may be reproduced or transmitted in any form or by any      //
//  means, electronic or mechanical, including photocopying, recording, or any   //
//  information storage and retrieval system in violation of the license under   //
//  which the source code is released.                                           //
//                                                                               //
//  The source code contained herein is free; it may be studied, copied,         //
// compiled and executed only for academic, non-commercial research purposes,    //
//  subject to the restrictions in YanSolutions License.                         //
//                                                                               //
//  You may not Re-distribute this VIP in any form for any purposes. Examples    //
//  of purposes would be running business operations, licensing,                 //
//  leasing, or selling the FreeVIP, distributing the FreeVIP for use            //
//  with commercial or non-commercial products, using the FreeVIP in             //
//  the creation or use of commercial or non-commercial products.                //
//                                                                               //
// THIS CODE IS PROVIDED ''AS IS'' AND WITHOUT ANY                               //
// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED                     //
// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A               //
// PARTICULAR PURPOSE. IN NO EVENT SHALL YS NOR ANY CONTRIBUTOR TO               //
// THE FREEVIP WILL BE LIABLE FOR ANY DAMAGES RELATED TO THE FREEVIP OR          //
// THIS LICENSE, INCLUDING DIRECT, INDIRECT, SPECIAL, CONSEQUENTIAL OR           //
// INCIDENTAL DAMAGES, TO THE MAXIMUM EXTENT THE LAW PERMITS, NO MATTER WHAT     //
// LEGAL THEORY IT IS BASED ON. ALSO, YOU MUST PASS THIS LIMITATION OF           //
// LIABILITY ON WHENEVER YOU DISTRIBUTE THE FREEVIP OR DERIVATIVE WORKS.         //
//                                                                               //
//  YanSolutions, Inc.                                                           //
//  Yerevan, Davidashen 4, 21/2                                                  //
//  Armenia, www.yansolutions.com                                                //
//                                                                               //
/////////////////////////////////////////////////////////////////////////////////// 

class seqItem extends uvm_sequence_item;
`uvm_object_utils(seqItem)

logic [8-1:0] rdata;
logic wfull;
logic rempty;
rand logic [8-1:0] wdata;
logic winc, wrst_n;
logic rinc, rrst_n;

fifoVerif_pkg::operation op;

function new (string name="seqItem");
	super.new(name);
endfunction


function void do_copy(uvm_object rhs);
		seqItem tr;
		if(!$cast(tr, rhs)) `uvm_fatal("trans1", "ILLEGAL do_copy() cast")
		rdata = tr.rdata;
		wfull = tr.wfull;
		rempty = tr.rempty;
		wdata = tr.wdata;
		winc = tr.winc;
		wrst_n = tr.wrst_n;
		rinc = tr.rinc;
		rrst_n = tr.rrst_n;
 endfunction 
 
  function bit do_compare(uvm_object rhs, uvm_comparer comparer= null);
		seqItem tr;
		bit eq;
		if(!$cast(tr, rhs)) `uvm_fatal("trans1", "ILLEGAL do_compare() cast")
		eq = super.do_compare(rhs, comparer);
		if (|rdata && |tr.rdata == "x")
				eq &= (rdata == tr.rdata);
		if (|wfull && |tr.wfull == "x")
				eq &= (wfull == tr.wfull);
		if (|wdata && |tr.wdata == "x")
				eq &= (wdata == tr.wdata);				
		if (|rempty && |tr.rempty == "x")
				eq &= (rempty == tr.rempty);
		return(eq);
 endfunction 
 
endclass