class writeFullSeq extends uvm_sequence #(seqItem);


endclass