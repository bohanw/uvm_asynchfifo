class writeTest extends uvm_test;
	`uvm_component_utils(writeTest)

	env env_h;



endclass
