module top();
	import uvm_pkg::*;


	`include "uvm_macros.svh";

	


endmodule // top